`define FREQ_INC_BITS 17
