`include "parameters.vh"
module SineLogTable(
    input  clk,
    input  [7:0] addr,
    output reg [9:0] value
);  

reg [9:0] sine_log_table[0:255];
initial begin
    sine_log_table[8'h000] <= 10'h3ff; sine_log_table[8'h001] <= 10'h33c; sine_log_table[8'h002] <= 10'h2e2; sine_log_table[8'h003] <= 10'h2a7; sine_log_table[8'h004] <= 10'h27a; sine_log_table[8'h005] <= 10'h257; sine_log_table[8'h006] <= 10'h239; sine_log_table[8'h007] <= 10'h220; sine_log_table[8'h008] <= 10'h20a; sine_log_table[8'h009] <= 10'h1f6; sine_log_table[8'h00a] <= 10'h1e4; sine_log_table[8'h00b] <= 10'h1d4; sine_log_table[8'h00c] <= 10'h1c6; sine_log_table[8'h00d] <= 10'h1b8; sine_log_table[8'h00e] <= 10'h1ab; sine_log_table[8'h00f] <= 10'h1a0;
    sine_log_table[8'h010] <= 10'h195; sine_log_table[8'h011] <= 10'h18a; sine_log_table[8'h012] <= 10'h181; sine_log_table[8'h013] <= 10'h177; sine_log_table[8'h014] <= 10'h16e; sine_log_table[8'h015] <= 10'h166; sine_log_table[8'h016] <= 10'h15e; sine_log_table[8'h017] <= 10'h156; sine_log_table[8'h018] <= 10'h14f; sine_log_table[8'h019] <= 10'h148; sine_log_table[8'h01a] <= 10'h141; sine_log_table[8'h01b] <= 10'h13b; sine_log_table[8'h01c] <= 10'h135; sine_log_table[8'h01d] <= 10'h12f; sine_log_table[8'h01e] <= 10'h129; sine_log_table[8'h01f] <= 10'h123;
    sine_log_table[8'h020] <= 10'h11e; sine_log_table[8'h021] <= 10'h118; sine_log_table[8'h022] <= 10'h113; sine_log_table[8'h023] <= 10'h10e; sine_log_table[8'h024] <= 10'h109; sine_log_table[8'h025] <= 10'h105; sine_log_table[8'h026] <= 10'h100; sine_log_table[8'h027] <= 10'h0fc; sine_log_table[8'h028] <= 10'h0f7; sine_log_table[8'h029] <= 10'h0f3; sine_log_table[8'h02a] <= 10'h0ef; sine_log_table[8'h02b] <= 10'h0eb; sine_log_table[8'h02c] <= 10'h0e7; sine_log_table[8'h02d] <= 10'h0e3; sine_log_table[8'h02e] <= 10'h0e0; sine_log_table[8'h02f] <= 10'h0dc;
    sine_log_table[8'h030] <= 10'h0d8; sine_log_table[8'h031] <= 10'h0d5; sine_log_table[8'h032] <= 10'h0d1; sine_log_table[8'h033] <= 10'h0ce; sine_log_table[8'h034] <= 10'h0cb; sine_log_table[8'h035] <= 10'h0c8; sine_log_table[8'h036] <= 10'h0c4; sine_log_table[8'h037] <= 10'h0c1; sine_log_table[8'h038] <= 10'h0be; sine_log_table[8'h039] <= 10'h0bb; sine_log_table[8'h03a] <= 10'h0b8; sine_log_table[8'h03b] <= 10'h0b6; sine_log_table[8'h03c] <= 10'h0b3; sine_log_table[8'h03d] <= 10'h0b0; sine_log_table[8'h03e] <= 10'h0ad; sine_log_table[8'h03f] <= 10'h0ab;
    sine_log_table[8'h040] <= 10'h0a8; sine_log_table[8'h041] <= 10'h0a5; sine_log_table[8'h042] <= 10'h0a3; sine_log_table[8'h043] <= 10'h0a0; sine_log_table[8'h044] <= 10'h09e; sine_log_table[8'h045] <= 10'h09c; sine_log_table[8'h046] <= 10'h099; sine_log_table[8'h047] <= 10'h097; sine_log_table[8'h048] <= 10'h095; sine_log_table[8'h049] <= 10'h092; sine_log_table[8'h04a] <= 10'h090; sine_log_table[8'h04b] <= 10'h08e; sine_log_table[8'h04c] <= 10'h08c; sine_log_table[8'h04d] <= 10'h08a; sine_log_table[8'h04e] <= 10'h088; sine_log_table[8'h04f] <= 10'h085;
    sine_log_table[8'h050] <= 10'h083; sine_log_table[8'h051] <= 10'h081; sine_log_table[8'h052] <= 10'h07f; sine_log_table[8'h053] <= 10'h07e; sine_log_table[8'h054] <= 10'h07c; sine_log_table[8'h055] <= 10'h07a; sine_log_table[8'h056] <= 10'h078; sine_log_table[8'h057] <= 10'h076; sine_log_table[8'h058] <= 10'h074; sine_log_table[8'h059] <= 10'h072; sine_log_table[8'h05a] <= 10'h071; sine_log_table[8'h05b] <= 10'h06f; sine_log_table[8'h05c] <= 10'h06d; sine_log_table[8'h05d] <= 10'h06c; sine_log_table[8'h05e] <= 10'h06a; sine_log_table[8'h05f] <= 10'h068;
    sine_log_table[8'h060] <= 10'h067; sine_log_table[8'h061] <= 10'h065; sine_log_table[8'h062] <= 10'h063; sine_log_table[8'h063] <= 10'h062; sine_log_table[8'h064] <= 10'h060; sine_log_table[8'h065] <= 10'h05f; sine_log_table[8'h066] <= 10'h05d; sine_log_table[8'h067] <= 10'h05c; sine_log_table[8'h068] <= 10'h05a; sine_log_table[8'h069] <= 10'h059; sine_log_table[8'h06a] <= 10'h057; sine_log_table[8'h06b] <= 10'h056; sine_log_table[8'h06c] <= 10'h055; sine_log_table[8'h06d] <= 10'h053; sine_log_table[8'h06e] <= 10'h052; sine_log_table[8'h06f] <= 10'h051;
    sine_log_table[8'h070] <= 10'h04f; sine_log_table[8'h071] <= 10'h04e; sine_log_table[8'h072] <= 10'h04d; sine_log_table[8'h073] <= 10'h04b; sine_log_table[8'h074] <= 10'h04a; sine_log_table[8'h075] <= 10'h049; sine_log_table[8'h076] <= 10'h048; sine_log_table[8'h077] <= 10'h046; sine_log_table[8'h078] <= 10'h045; sine_log_table[8'h079] <= 10'h044; sine_log_table[8'h07a] <= 10'h043; sine_log_table[8'h07b] <= 10'h042; sine_log_table[8'h07c] <= 10'h041; sine_log_table[8'h07d] <= 10'h040; sine_log_table[8'h07e] <= 10'h03e; sine_log_table[8'h07f] <= 10'h03d;
    sine_log_table[8'h080] <= 10'h03c; sine_log_table[8'h081] <= 10'h03b; sine_log_table[8'h082] <= 10'h03a; sine_log_table[8'h083] <= 10'h039; sine_log_table[8'h084] <= 10'h038; sine_log_table[8'h085] <= 10'h037; sine_log_table[8'h086] <= 10'h036; sine_log_table[8'h087] <= 10'h035; sine_log_table[8'h088] <= 10'h034; sine_log_table[8'h089] <= 10'h033; sine_log_table[8'h08a] <= 10'h032; sine_log_table[8'h08b] <= 10'h031; sine_log_table[8'h08c] <= 10'h030; sine_log_table[8'h08d] <= 10'h02f; sine_log_table[8'h08e] <= 10'h02e; sine_log_table[8'h08f] <= 10'h02d;
    sine_log_table[8'h090] <= 10'h02d; sine_log_table[8'h091] <= 10'h02c; sine_log_table[8'h092] <= 10'h02b; sine_log_table[8'h093] <= 10'h02a; sine_log_table[8'h094] <= 10'h029; sine_log_table[8'h095] <= 10'h028; sine_log_table[8'h096] <= 10'h027; sine_log_table[8'h097] <= 10'h027; sine_log_table[8'h098] <= 10'h026; sine_log_table[8'h099] <= 10'h025; sine_log_table[8'h09a] <= 10'h024; sine_log_table[8'h09b] <= 10'h023; sine_log_table[8'h09c] <= 10'h023; sine_log_table[8'h09d] <= 10'h022; sine_log_table[8'h09e] <= 10'h021; sine_log_table[8'h09f] <= 10'h020;
    sine_log_table[8'h0a0] <= 10'h020; sine_log_table[8'h0a1] <= 10'h01f; sine_log_table[8'h0a2] <= 10'h01e; sine_log_table[8'h0a3] <= 10'h01e; sine_log_table[8'h0a4] <= 10'h01d; sine_log_table[8'h0a5] <= 10'h01c; sine_log_table[8'h0a6] <= 10'h01c; sine_log_table[8'h0a7] <= 10'h01b; sine_log_table[8'h0a8] <= 10'h01a; sine_log_table[8'h0a9] <= 10'h01a; sine_log_table[8'h0aa] <= 10'h019; sine_log_table[8'h0ab] <= 10'h018; sine_log_table[8'h0ac] <= 10'h018; sine_log_table[8'h0ad] <= 10'h017; sine_log_table[8'h0ae] <= 10'h017; sine_log_table[8'h0af] <= 10'h016;
    sine_log_table[8'h0b0] <= 10'h015; sine_log_table[8'h0b1] <= 10'h015; sine_log_table[8'h0b2] <= 10'h014; sine_log_table[8'h0b3] <= 10'h014; sine_log_table[8'h0b4] <= 10'h013; sine_log_table[8'h0b5] <= 10'h013; sine_log_table[8'h0b6] <= 10'h012; sine_log_table[8'h0b7] <= 10'h012; sine_log_table[8'h0b8] <= 10'h011; sine_log_table[8'h0b9] <= 10'h011; sine_log_table[8'h0ba] <= 10'h010; sine_log_table[8'h0bb] <= 10'h010; sine_log_table[8'h0bc] <= 10'h00f; sine_log_table[8'h0bd] <= 10'h00f; sine_log_table[8'h0be] <= 10'h00e; sine_log_table[8'h0bf] <= 10'h00e;
    sine_log_table[8'h0c0] <= 10'h00d; sine_log_table[8'h0c1] <= 10'h00d; sine_log_table[8'h0c2] <= 10'h00c; sine_log_table[8'h0c3] <= 10'h00c; sine_log_table[8'h0c4] <= 10'h00c; sine_log_table[8'h0c5] <= 10'h00b; sine_log_table[8'h0c6] <= 10'h00b; sine_log_table[8'h0c7] <= 10'h00a; sine_log_table[8'h0c8] <= 10'h00a; sine_log_table[8'h0c9] <= 10'h00a; sine_log_table[8'h0ca] <= 10'h009; sine_log_table[8'h0cb] <= 10'h009; sine_log_table[8'h0cc] <= 10'h008; sine_log_table[8'h0cd] <= 10'h008; sine_log_table[8'h0ce] <= 10'h008; sine_log_table[8'h0cf] <= 10'h007;
    sine_log_table[8'h0d0] <= 10'h007; sine_log_table[8'h0d1] <= 10'h007; sine_log_table[8'h0d2] <= 10'h006; sine_log_table[8'h0d3] <= 10'h006; sine_log_table[8'h0d4] <= 10'h006; sine_log_table[8'h0d5] <= 10'h006; sine_log_table[8'h0d6] <= 10'h005; sine_log_table[8'h0d7] <= 10'h005; sine_log_table[8'h0d8] <= 10'h005; sine_log_table[8'h0d9] <= 10'h004; sine_log_table[8'h0da] <= 10'h004; sine_log_table[8'h0db] <= 10'h004; sine_log_table[8'h0dc] <= 10'h004; sine_log_table[8'h0dd] <= 10'h003; sine_log_table[8'h0de] <= 10'h003; sine_log_table[8'h0df] <= 10'h003;
    sine_log_table[8'h0e0] <= 10'h003; sine_log_table[8'h0e1] <= 10'h003; sine_log_table[8'h0e2] <= 10'h002; sine_log_table[8'h0e3] <= 10'h002; sine_log_table[8'h0e4] <= 10'h002; sine_log_table[8'h0e5] <= 10'h002; sine_log_table[8'h0e6] <= 10'h002; sine_log_table[8'h0e7] <= 10'h002; sine_log_table[8'h0e8] <= 10'h001; sine_log_table[8'h0e9] <= 10'h001; sine_log_table[8'h0ea] <= 10'h001; sine_log_table[8'h0eb] <= 10'h001; sine_log_table[8'h0ec] <= 10'h001; sine_log_table[8'h0ed] <= 10'h001; sine_log_table[8'h0ee] <= 10'h001; sine_log_table[8'h0ef] <= 10'h000;
    sine_log_table[8'h0f0] <= 10'h000; sine_log_table[8'h0f1] <= 10'h000; sine_log_table[8'h0f2] <= 10'h000; sine_log_table[8'h0f3] <= 10'h000; sine_log_table[8'h0f4] <= 10'h000; sine_log_table[8'h0f5] <= 10'h000; sine_log_table[8'h0f6] <= 10'h000; sine_log_table[8'h0f7] <= 10'h000; sine_log_table[8'h0f8] <= 10'h000; sine_log_table[8'h0f9] <= 10'h000; sine_log_table[8'h0fa] <= 10'h000; sine_log_table[8'h0fb] <= 10'h000; sine_log_table[8'h0fc] <= 10'h000; sine_log_table[8'h0fd] <= 10'h000; sine_log_table[8'h0fe] <= 10'h000; sine_log_table[8'h0ff] <= 10'h000;
end

always @ (posedge clk) begin
    value <= sine_log_table[addr];
end

endmodule

module ExpTable(
    input  clk,
    input  [11:0] addr,
    output reg [8:0] value
);  

reg [8:0] exp_table[0:1535];
initial begin
    exp_table[11'h000] <= 9'h1ff; exp_table[11'h001] <= 9'h1fc; exp_table[11'h002] <= 9'h1f9; exp_table[11'h003] <= 9'h1f6; exp_table[11'h004] <= 9'h1f3; exp_table[11'h005] <= 9'h1f0; exp_table[11'h006] <= 9'h1ed; exp_table[11'h007] <= 9'h1eb; exp_table[11'h008] <= 9'h1e8; exp_table[11'h009] <= 9'h1e5; exp_table[11'h00a] <= 9'h1e2; exp_table[11'h00b] <= 9'h1e0; exp_table[11'h00c] <= 9'h1dd; exp_table[11'h00d] <= 9'h1da; exp_table[11'h00e] <= 9'h1d8; exp_table[11'h00f] <= 9'h1d5;
    exp_table[11'h010] <= 9'h1d2; exp_table[11'h011] <= 9'h1d0; exp_table[11'h012] <= 9'h1cd; exp_table[11'h013] <= 9'h1ca; exp_table[11'h014] <= 9'h1c8; exp_table[11'h015] <= 9'h1c5; exp_table[11'h016] <= 9'h1c3; exp_table[11'h017] <= 9'h1c0; exp_table[11'h018] <= 9'h1be; exp_table[11'h019] <= 9'h1bb; exp_table[11'h01a] <= 9'h1b9; exp_table[11'h01b] <= 9'h1b6; exp_table[11'h01c] <= 9'h1b4; exp_table[11'h01d] <= 9'h1b1; exp_table[11'h01e] <= 9'h1af; exp_table[11'h01f] <= 9'h1ac;
    exp_table[11'h020] <= 9'h1aa; exp_table[11'h021] <= 9'h1a7; exp_table[11'h022] <= 9'h1a5; exp_table[11'h023] <= 9'h1a3; exp_table[11'h024] <= 9'h1a0; exp_table[11'h025] <= 9'h19e; exp_table[11'h026] <= 9'h19c; exp_table[11'h027] <= 9'h199; exp_table[11'h028] <= 9'h197; exp_table[11'h029] <= 9'h195; exp_table[11'h02a] <= 9'h192; exp_table[11'h02b] <= 9'h190; exp_table[11'h02c] <= 9'h18e; exp_table[11'h02d] <= 9'h18c; exp_table[11'h02e] <= 9'h189; exp_table[11'h02f] <= 9'h187;
    exp_table[11'h030] <= 9'h185; exp_table[11'h031] <= 9'h183; exp_table[11'h032] <= 9'h181; exp_table[11'h033] <= 9'h17e; exp_table[11'h034] <= 9'h17c; exp_table[11'h035] <= 9'h17a; exp_table[11'h036] <= 9'h178; exp_table[11'h037] <= 9'h176; exp_table[11'h038] <= 9'h174; exp_table[11'h039] <= 9'h172; exp_table[11'h03a] <= 9'h170; exp_table[11'h03b] <= 9'h16d; exp_table[11'h03c] <= 9'h16b; exp_table[11'h03d] <= 9'h169; exp_table[11'h03e] <= 9'h167; exp_table[11'h03f] <= 9'h165;
    exp_table[11'h040] <= 9'h163; exp_table[11'h041] <= 9'h161; exp_table[11'h042] <= 9'h15f; exp_table[11'h043] <= 9'h15d; exp_table[11'h044] <= 9'h15b; exp_table[11'h045] <= 9'h159; exp_table[11'h046] <= 9'h157; exp_table[11'h047] <= 9'h155; exp_table[11'h048] <= 9'h154; exp_table[11'h049] <= 9'h152; exp_table[11'h04a] <= 9'h150; exp_table[11'h04b] <= 9'h14e; exp_table[11'h04c] <= 9'h14c; exp_table[11'h04d] <= 9'h14a; exp_table[11'h04e] <= 9'h148; exp_table[11'h04f] <= 9'h146;
    exp_table[11'h050] <= 9'h145; exp_table[11'h051] <= 9'h143; exp_table[11'h052] <= 9'h141; exp_table[11'h053] <= 9'h13f; exp_table[11'h054] <= 9'h13d; exp_table[11'h055] <= 9'h13b; exp_table[11'h056] <= 9'h13a; exp_table[11'h057] <= 9'h138; exp_table[11'h058] <= 9'h136; exp_table[11'h059] <= 9'h134; exp_table[11'h05a] <= 9'h133; exp_table[11'h05b] <= 9'h131; exp_table[11'h05c] <= 9'h12f; exp_table[11'h05d] <= 9'h12d; exp_table[11'h05e] <= 9'h12c; exp_table[11'h05f] <= 9'h12a;
    exp_table[11'h060] <= 9'h128; exp_table[11'h061] <= 9'h127; exp_table[11'h062] <= 9'h125; exp_table[11'h063] <= 9'h123; exp_table[11'h064] <= 9'h122; exp_table[11'h065] <= 9'h120; exp_table[11'h066] <= 9'h11e; exp_table[11'h067] <= 9'h11d; exp_table[11'h068] <= 9'h11b; exp_table[11'h069] <= 9'h11a; exp_table[11'h06a] <= 9'h118; exp_table[11'h06b] <= 9'h116; exp_table[11'h06c] <= 9'h115; exp_table[11'h06d] <= 9'h113; exp_table[11'h06e] <= 9'h112; exp_table[11'h06f] <= 9'h110;
    exp_table[11'h070] <= 9'h10f; exp_table[11'h071] <= 9'h10d; exp_table[11'h072] <= 9'h10c; exp_table[11'h073] <= 9'h10a; exp_table[11'h074] <= 9'h109; exp_table[11'h075] <= 9'h107; exp_table[11'h076] <= 9'h106; exp_table[11'h077] <= 9'h104; exp_table[11'h078] <= 9'h103; exp_table[11'h079] <= 9'h101; exp_table[11'h07a] <= 9'h100; exp_table[11'h07b] <= 9'h0fe; exp_table[11'h07c] <= 9'h0fd; exp_table[11'h07d] <= 9'h0fb; exp_table[11'h07e] <= 9'h0fa; exp_table[11'h07f] <= 9'h0f9;
    exp_table[11'h080] <= 9'h0f7; exp_table[11'h081] <= 9'h0f6; exp_table[11'h082] <= 9'h0f4; exp_table[11'h083] <= 9'h0f3; exp_table[11'h084] <= 9'h0f2; exp_table[11'h085] <= 9'h0f0; exp_table[11'h086] <= 9'h0ef; exp_table[11'h087] <= 9'h0ee; exp_table[11'h088] <= 9'h0ec; exp_table[11'h089] <= 9'h0eb; exp_table[11'h08a] <= 9'h0ea; exp_table[11'h08b] <= 9'h0e8; exp_table[11'h08c] <= 9'h0e7; exp_table[11'h08d] <= 9'h0e6; exp_table[11'h08e] <= 9'h0e4; exp_table[11'h08f] <= 9'h0e3;
    exp_table[11'h090] <= 9'h0e2; exp_table[11'h091] <= 9'h0e1; exp_table[11'h092] <= 9'h0df; exp_table[11'h093] <= 9'h0de; exp_table[11'h094] <= 9'h0dd; exp_table[11'h095] <= 9'h0db; exp_table[11'h096] <= 9'h0da; exp_table[11'h097] <= 9'h0d9; exp_table[11'h098] <= 9'h0d8; exp_table[11'h099] <= 9'h0d7; exp_table[11'h09a] <= 9'h0d5; exp_table[11'h09b] <= 9'h0d4; exp_table[11'h09c] <= 9'h0d3; exp_table[11'h09d] <= 9'h0d2; exp_table[11'h09e] <= 9'h0d1; exp_table[11'h09f] <= 9'h0cf;
    exp_table[11'h0a0] <= 9'h0ce; exp_table[11'h0a1] <= 9'h0cd; exp_table[11'h0a2] <= 9'h0cc; exp_table[11'h0a3] <= 9'h0cb; exp_table[11'h0a4] <= 9'h0ca; exp_table[11'h0a5] <= 9'h0c8; exp_table[11'h0a6] <= 9'h0c7; exp_table[11'h0a7] <= 9'h0c6; exp_table[11'h0a8] <= 9'h0c5; exp_table[11'h0a9] <= 9'h0c4; exp_table[11'h0aa] <= 9'h0c3; exp_table[11'h0ab] <= 9'h0c2; exp_table[11'h0ac] <= 9'h0c1; exp_table[11'h0ad] <= 9'h0c0; exp_table[11'h0ae] <= 9'h0be; exp_table[11'h0af] <= 9'h0bd;
    exp_table[11'h0b0] <= 9'h0bc; exp_table[11'h0b1] <= 9'h0bb; exp_table[11'h0b2] <= 9'h0ba; exp_table[11'h0b3] <= 9'h0b9; exp_table[11'h0b4] <= 9'h0b8; exp_table[11'h0b5] <= 9'h0b7; exp_table[11'h0b6] <= 9'h0b6; exp_table[11'h0b7] <= 9'h0b5; exp_table[11'h0b8] <= 9'h0b4; exp_table[11'h0b9] <= 9'h0b3; exp_table[11'h0ba] <= 9'h0b2; exp_table[11'h0bb] <= 9'h0b1; exp_table[11'h0bc] <= 9'h0b0; exp_table[11'h0bd] <= 9'h0af; exp_table[11'h0be] <= 9'h0ae; exp_table[11'h0bf] <= 9'h0ad;
    exp_table[11'h0c0] <= 9'h0ac; exp_table[11'h0c1] <= 9'h0ab; exp_table[11'h0c2] <= 9'h0aa; exp_table[11'h0c3] <= 9'h0a9; exp_table[11'h0c4] <= 9'h0a8; exp_table[11'h0c5] <= 9'h0a7; exp_table[11'h0c6] <= 9'h0a6; exp_table[11'h0c7] <= 9'h0a5; exp_table[11'h0c8] <= 9'h0a4; exp_table[11'h0c9] <= 9'h0a3; exp_table[11'h0ca] <= 9'h0a2; exp_table[11'h0cb] <= 9'h0a2; exp_table[11'h0cc] <= 9'h0a1; exp_table[11'h0cd] <= 9'h0a0; exp_table[11'h0ce] <= 9'h09f; exp_table[11'h0cf] <= 9'h09e;
    exp_table[11'h0d0] <= 9'h09d; exp_table[11'h0d1] <= 9'h09c; exp_table[11'h0d2] <= 9'h09b; exp_table[11'h0d3] <= 9'h09a; exp_table[11'h0d4] <= 9'h09a; exp_table[11'h0d5] <= 9'h099; exp_table[11'h0d6] <= 9'h098; exp_table[11'h0d7] <= 9'h097; exp_table[11'h0d8] <= 9'h096; exp_table[11'h0d9] <= 9'h095; exp_table[11'h0da] <= 9'h094; exp_table[11'h0db] <= 9'h094; exp_table[11'h0dc] <= 9'h093; exp_table[11'h0dd] <= 9'h092; exp_table[11'h0de] <= 9'h091; exp_table[11'h0df] <= 9'h090;
    exp_table[11'h0e0] <= 9'h08f; exp_table[11'h0e1] <= 9'h08f; exp_table[11'h0e2] <= 9'h08e; exp_table[11'h0e3] <= 9'h08d; exp_table[11'h0e4] <= 9'h08c; exp_table[11'h0e5] <= 9'h08b; exp_table[11'h0e6] <= 9'h08b; exp_table[11'h0e7] <= 9'h08a; exp_table[11'h0e8] <= 9'h089; exp_table[11'h0e9] <= 9'h088; exp_table[11'h0ea] <= 9'h088; exp_table[11'h0eb] <= 9'h087; exp_table[11'h0ec] <= 9'h086; exp_table[11'h0ed] <= 9'h085; exp_table[11'h0ee] <= 9'h084; exp_table[11'h0ef] <= 9'h084;
    exp_table[11'h0f0] <= 9'h083; exp_table[11'h0f1] <= 9'h082; exp_table[11'h0f2] <= 9'h081; exp_table[11'h0f3] <= 9'h081; exp_table[11'h0f4] <= 9'h080; exp_table[11'h0f5] <= 9'h07f; exp_table[11'h0f6] <= 9'h07f; exp_table[11'h0f7] <= 9'h07e; exp_table[11'h0f8] <= 9'h07d; exp_table[11'h0f9] <= 9'h07c; exp_table[11'h0fa] <= 9'h07c; exp_table[11'h0fb] <= 9'h07b; exp_table[11'h0fc] <= 9'h07a; exp_table[11'h0fd] <= 9'h07a; exp_table[11'h0fe] <= 9'h079; exp_table[11'h0ff] <= 9'h078;
    exp_table[11'h100] <= 9'h078; exp_table[11'h101] <= 9'h077; exp_table[11'h102] <= 9'h076; exp_table[11'h103] <= 9'h076; exp_table[11'h104] <= 9'h075; exp_table[11'h105] <= 9'h074; exp_table[11'h106] <= 9'h074; exp_table[11'h107] <= 9'h073; exp_table[11'h108] <= 9'h072; exp_table[11'h109] <= 9'h072; exp_table[11'h10a] <= 9'h071; exp_table[11'h10b] <= 9'h070; exp_table[11'h10c] <= 9'h070; exp_table[11'h10d] <= 9'h06f; exp_table[11'h10e] <= 9'h06e; exp_table[11'h10f] <= 9'h06e;
    exp_table[11'h110] <= 9'h06d; exp_table[11'h111] <= 9'h06d; exp_table[11'h112] <= 9'h06c; exp_table[11'h113] <= 9'h06b; exp_table[11'h114] <= 9'h06b; exp_table[11'h115] <= 9'h06a; exp_table[11'h116] <= 9'h06a; exp_table[11'h117] <= 9'h069; exp_table[11'h118] <= 9'h068; exp_table[11'h119] <= 9'h068; exp_table[11'h11a] <= 9'h067; exp_table[11'h11b] <= 9'h067; exp_table[11'h11c] <= 9'h066; exp_table[11'h11d] <= 9'h065; exp_table[11'h11e] <= 9'h065; exp_table[11'h11f] <= 9'h064;
    exp_table[11'h120] <= 9'h064; exp_table[11'h121] <= 9'h063; exp_table[11'h122] <= 9'h063; exp_table[11'h123] <= 9'h062; exp_table[11'h124] <= 9'h061; exp_table[11'h125] <= 9'h061; exp_table[11'h126] <= 9'h060; exp_table[11'h127] <= 9'h060; exp_table[11'h128] <= 9'h05f; exp_table[11'h129] <= 9'h05f; exp_table[11'h12a] <= 9'h05e; exp_table[11'h12b] <= 9'h05e; exp_table[11'h12c] <= 9'h05d; exp_table[11'h12d] <= 9'h05d; exp_table[11'h12e] <= 9'h05c; exp_table[11'h12f] <= 9'h05c;
    exp_table[11'h130] <= 9'h05b; exp_table[11'h131] <= 9'h05b; exp_table[11'h132] <= 9'h05a; exp_table[11'h133] <= 9'h059; exp_table[11'h134] <= 9'h059; exp_table[11'h135] <= 9'h058; exp_table[11'h136] <= 9'h058; exp_table[11'h137] <= 9'h057; exp_table[11'h138] <= 9'h057; exp_table[11'h139] <= 9'h056; exp_table[11'h13a] <= 9'h056; exp_table[11'h13b] <= 9'h056; exp_table[11'h13c] <= 9'h055; exp_table[11'h13d] <= 9'h055; exp_table[11'h13e] <= 9'h054; exp_table[11'h13f] <= 9'h054;
    exp_table[11'h140] <= 9'h053; exp_table[11'h141] <= 9'h053; exp_table[11'h142] <= 9'h052; exp_table[11'h143] <= 9'h052; exp_table[11'h144] <= 9'h051; exp_table[11'h145] <= 9'h051; exp_table[11'h146] <= 9'h050; exp_table[11'h147] <= 9'h050; exp_table[11'h148] <= 9'h04f; exp_table[11'h149] <= 9'h04f; exp_table[11'h14a] <= 9'h04f; exp_table[11'h14b] <= 9'h04e; exp_table[11'h14c] <= 9'h04e; exp_table[11'h14d] <= 9'h04d; exp_table[11'h14e] <= 9'h04d; exp_table[11'h14f] <= 9'h04c;
    exp_table[11'h150] <= 9'h04c; exp_table[11'h151] <= 9'h04b; exp_table[11'h152] <= 9'h04b; exp_table[11'h153] <= 9'h04b; exp_table[11'h154] <= 9'h04a; exp_table[11'h155] <= 9'h04a; exp_table[11'h156] <= 9'h049; exp_table[11'h157] <= 9'h049; exp_table[11'h158] <= 9'h049; exp_table[11'h159] <= 9'h048; exp_table[11'h15a] <= 9'h048; exp_table[11'h15b] <= 9'h047; exp_table[11'h15c] <= 9'h047; exp_table[11'h15d] <= 9'h046; exp_table[11'h15e] <= 9'h046; exp_table[11'h15f] <= 9'h046;
    exp_table[11'h160] <= 9'h045; exp_table[11'h161] <= 9'h045; exp_table[11'h162] <= 9'h044; exp_table[11'h163] <= 9'h044; exp_table[11'h164] <= 9'h044; exp_table[11'h165] <= 9'h043; exp_table[11'h166] <= 9'h043; exp_table[11'h167] <= 9'h043; exp_table[11'h168] <= 9'h042; exp_table[11'h169] <= 9'h042; exp_table[11'h16a] <= 9'h041; exp_table[11'h16b] <= 9'h041; exp_table[11'h16c] <= 9'h041; exp_table[11'h16d] <= 9'h040; exp_table[11'h16e] <= 9'h040; exp_table[11'h16f] <= 9'h040;
    exp_table[11'h170] <= 9'h03f; exp_table[11'h171] <= 9'h03f; exp_table[11'h172] <= 9'h03f; exp_table[11'h173] <= 9'h03e; exp_table[11'h174] <= 9'h03e; exp_table[11'h175] <= 9'h03d; exp_table[11'h176] <= 9'h03d; exp_table[11'h177] <= 9'h03d; exp_table[11'h178] <= 9'h03c; exp_table[11'h179] <= 9'h03c; exp_table[11'h17a] <= 9'h03c; exp_table[11'h17b] <= 9'h03b; exp_table[11'h17c] <= 9'h03b; exp_table[11'h17d] <= 9'h03b; exp_table[11'h17e] <= 9'h03a; exp_table[11'h17f] <= 9'h03a;
    exp_table[11'h180] <= 9'h03a; exp_table[11'h181] <= 9'h039; exp_table[11'h182] <= 9'h039; exp_table[11'h183] <= 9'h039; exp_table[11'h184] <= 9'h038; exp_table[11'h185] <= 9'h038; exp_table[11'h186] <= 9'h038; exp_table[11'h187] <= 9'h037; exp_table[11'h188] <= 9'h037; exp_table[11'h189] <= 9'h037; exp_table[11'h18a] <= 9'h037; exp_table[11'h18b] <= 9'h036; exp_table[11'h18c] <= 9'h036; exp_table[11'h18d] <= 9'h036; exp_table[11'h18e] <= 9'h035; exp_table[11'h18f] <= 9'h035;
    exp_table[11'h190] <= 9'h035; exp_table[11'h191] <= 9'h034; exp_table[11'h192] <= 9'h034; exp_table[11'h193] <= 9'h034; exp_table[11'h194] <= 9'h033; exp_table[11'h195] <= 9'h033; exp_table[11'h196] <= 9'h033; exp_table[11'h197] <= 9'h033; exp_table[11'h198] <= 9'h032; exp_table[11'h199] <= 9'h032; exp_table[11'h19a] <= 9'h032; exp_table[11'h19b] <= 9'h031; exp_table[11'h19c] <= 9'h031; exp_table[11'h19d] <= 9'h031; exp_table[11'h19e] <= 9'h031; exp_table[11'h19f] <= 9'h030;
    exp_table[11'h1a0] <= 9'h030; exp_table[11'h1a1] <= 9'h030; exp_table[11'h1a2] <= 9'h030; exp_table[11'h1a3] <= 9'h02f; exp_table[11'h1a4] <= 9'h02f; exp_table[11'h1a5] <= 9'h02f; exp_table[11'h1a6] <= 9'h02e; exp_table[11'h1a7] <= 9'h02e; exp_table[11'h1a8] <= 9'h02e; exp_table[11'h1a9] <= 9'h02e; exp_table[11'h1aa] <= 9'h02d; exp_table[11'h1ab] <= 9'h02d; exp_table[11'h1ac] <= 9'h02d; exp_table[11'h1ad] <= 9'h02d; exp_table[11'h1ae] <= 9'h02c; exp_table[11'h1af] <= 9'h02c;
    exp_table[11'h1b0] <= 9'h02c; exp_table[11'h1b1] <= 9'h02c; exp_table[11'h1b2] <= 9'h02b; exp_table[11'h1b3] <= 9'h02b; exp_table[11'h1b4] <= 9'h02b; exp_table[11'h1b5] <= 9'h02b; exp_table[11'h1b6] <= 9'h02a; exp_table[11'h1b7] <= 9'h02a; exp_table[11'h1b8] <= 9'h02a; exp_table[11'h1b9] <= 9'h02a; exp_table[11'h1ba] <= 9'h029; exp_table[11'h1bb] <= 9'h029; exp_table[11'h1bc] <= 9'h029; exp_table[11'h1bd] <= 9'h029; exp_table[11'h1be] <= 9'h028; exp_table[11'h1bf] <= 9'h028;
    exp_table[11'h1c0] <= 9'h028; exp_table[11'h1c1] <= 9'h028; exp_table[11'h1c2] <= 9'h028; exp_table[11'h1c3] <= 9'h027; exp_table[11'h1c4] <= 9'h027; exp_table[11'h1c5] <= 9'h027; exp_table[11'h1c6] <= 9'h027; exp_table[11'h1c7] <= 9'h026; exp_table[11'h1c8] <= 9'h026; exp_table[11'h1c9] <= 9'h026; exp_table[11'h1ca] <= 9'h026; exp_table[11'h1cb] <= 9'h026; exp_table[11'h1cc] <= 9'h025; exp_table[11'h1cd] <= 9'h025; exp_table[11'h1ce] <= 9'h025; exp_table[11'h1cf] <= 9'h025;
    exp_table[11'h1d0] <= 9'h025; exp_table[11'h1d1] <= 9'h024; exp_table[11'h1d2] <= 9'h024; exp_table[11'h1d3] <= 9'h024; exp_table[11'h1d4] <= 9'h024; exp_table[11'h1d5] <= 9'h023; exp_table[11'h1d6] <= 9'h023; exp_table[11'h1d7] <= 9'h023; exp_table[11'h1d8] <= 9'h023; exp_table[11'h1d9] <= 9'h023; exp_table[11'h1da] <= 9'h022; exp_table[11'h1db] <= 9'h022; exp_table[11'h1dc] <= 9'h022; exp_table[11'h1dd] <= 9'h022; exp_table[11'h1de] <= 9'h022; exp_table[11'h1df] <= 9'h022;
    exp_table[11'h1e0] <= 9'h021; exp_table[11'h1e1] <= 9'h021; exp_table[11'h1e2] <= 9'h021; exp_table[11'h1e3] <= 9'h021; exp_table[11'h1e4] <= 9'h021; exp_table[11'h1e5] <= 9'h020; exp_table[11'h1e6] <= 9'h020; exp_table[11'h1e7] <= 9'h020; exp_table[11'h1e8] <= 9'h020; exp_table[11'h1e9] <= 9'h020; exp_table[11'h1ea] <= 9'h01f; exp_table[11'h1eb] <= 9'h01f; exp_table[11'h1ec] <= 9'h01f; exp_table[11'h1ed] <= 9'h01f; exp_table[11'h1ee] <= 9'h01f; exp_table[11'h1ef] <= 9'h01f;
    exp_table[11'h1f0] <= 9'h01e; exp_table[11'h1f1] <= 9'h01e; exp_table[11'h1f2] <= 9'h01e; exp_table[11'h1f3] <= 9'h01e; exp_table[11'h1f4] <= 9'h01e; exp_table[11'h1f5] <= 9'h01e; exp_table[11'h1f6] <= 9'h01d; exp_table[11'h1f7] <= 9'h01d; exp_table[11'h1f8] <= 9'h01d; exp_table[11'h1f9] <= 9'h01d; exp_table[11'h1fa] <= 9'h01d; exp_table[11'h1fb] <= 9'h01d; exp_table[11'h1fc] <= 9'h01c; exp_table[11'h1fd] <= 9'h01c; exp_table[11'h1fe] <= 9'h01c; exp_table[11'h1ff] <= 9'h01c;
    exp_table[11'h200] <= 9'h01c; exp_table[11'h201] <= 9'h01c; exp_table[11'h202] <= 9'h01b; exp_table[11'h203] <= 9'h01b; exp_table[11'h204] <= 9'h01b; exp_table[11'h205] <= 9'h01b; exp_table[11'h206] <= 9'h01b; exp_table[11'h207] <= 9'h01b; exp_table[11'h208] <= 9'h01a; exp_table[11'h209] <= 9'h01a; exp_table[11'h20a] <= 9'h01a; exp_table[11'h20b] <= 9'h01a; exp_table[11'h20c] <= 9'h01a; exp_table[11'h20d] <= 9'h01a; exp_table[11'h20e] <= 9'h01a; exp_table[11'h20f] <= 9'h019;
    exp_table[11'h210] <= 9'h019; exp_table[11'h211] <= 9'h019; exp_table[11'h212] <= 9'h019; exp_table[11'h213] <= 9'h019; exp_table[11'h214] <= 9'h019; exp_table[11'h215] <= 9'h019; exp_table[11'h216] <= 9'h018; exp_table[11'h217] <= 9'h018; exp_table[11'h218] <= 9'h018; exp_table[11'h219] <= 9'h018; exp_table[11'h21a] <= 9'h018; exp_table[11'h21b] <= 9'h018; exp_table[11'h21c] <= 9'h018; exp_table[11'h21d] <= 9'h017; exp_table[11'h21e] <= 9'h017; exp_table[11'h21f] <= 9'h017;
    exp_table[11'h220] <= 9'h017; exp_table[11'h221] <= 9'h017; exp_table[11'h222] <= 9'h017; exp_table[11'h223] <= 9'h017; exp_table[11'h224] <= 9'h017; exp_table[11'h225] <= 9'h016; exp_table[11'h226] <= 9'h016; exp_table[11'h227] <= 9'h016; exp_table[11'h228] <= 9'h016; exp_table[11'h229] <= 9'h016; exp_table[11'h22a] <= 9'h016; exp_table[11'h22b] <= 9'h016; exp_table[11'h22c] <= 9'h016; exp_table[11'h22d] <= 9'h015; exp_table[11'h22e] <= 9'h015; exp_table[11'h22f] <= 9'h015;
    exp_table[11'h230] <= 9'h015; exp_table[11'h231] <= 9'h015; exp_table[11'h232] <= 9'h015; exp_table[11'h233] <= 9'h015; exp_table[11'h234] <= 9'h015; exp_table[11'h235] <= 9'h014; exp_table[11'h236] <= 9'h014; exp_table[11'h237] <= 9'h014; exp_table[11'h238] <= 9'h014; exp_table[11'h239] <= 9'h014; exp_table[11'h23a] <= 9'h014; exp_table[11'h23b] <= 9'h014; exp_table[11'h23c] <= 9'h014; exp_table[11'h23d] <= 9'h013; exp_table[11'h23e] <= 9'h013; exp_table[11'h23f] <= 9'h013;
    exp_table[11'h240] <= 9'h013; exp_table[11'h241] <= 9'h013; exp_table[11'h242] <= 9'h013; exp_table[11'h243] <= 9'h013; exp_table[11'h244] <= 9'h013; exp_table[11'h245] <= 9'h013; exp_table[11'h246] <= 9'h012; exp_table[11'h247] <= 9'h012; exp_table[11'h248] <= 9'h012; exp_table[11'h249] <= 9'h012; exp_table[11'h24a] <= 9'h012; exp_table[11'h24b] <= 9'h012; exp_table[11'h24c] <= 9'h012; exp_table[11'h24d] <= 9'h012; exp_table[11'h24e] <= 9'h012; exp_table[11'h24f] <= 9'h012;
    exp_table[11'h250] <= 9'h011; exp_table[11'h251] <= 9'h011; exp_table[11'h252] <= 9'h011; exp_table[11'h253] <= 9'h011; exp_table[11'h254] <= 9'h011; exp_table[11'h255] <= 9'h011; exp_table[11'h256] <= 9'h011; exp_table[11'h257] <= 9'h011; exp_table[11'h258] <= 9'h011; exp_table[11'h259] <= 9'h011; exp_table[11'h25a] <= 9'h010; exp_table[11'h25b] <= 9'h010; exp_table[11'h25c] <= 9'h010; exp_table[11'h25d] <= 9'h010; exp_table[11'h25e] <= 9'h010; exp_table[11'h25f] <= 9'h010;
    exp_table[11'h260] <= 9'h010; exp_table[11'h261] <= 9'h010; exp_table[11'h262] <= 9'h010; exp_table[11'h263] <= 9'h010; exp_table[11'h264] <= 9'h010; exp_table[11'h265] <= 9'h00f; exp_table[11'h266] <= 9'h00f; exp_table[11'h267] <= 9'h00f; exp_table[11'h268] <= 9'h00f; exp_table[11'h269] <= 9'h00f; exp_table[11'h26a] <= 9'h00f; exp_table[11'h26b] <= 9'h00f; exp_table[11'h26c] <= 9'h00f; exp_table[11'h26d] <= 9'h00f; exp_table[11'h26e] <= 9'h00f; exp_table[11'h26f] <= 9'h00f;
    exp_table[11'h270] <= 9'h00e; exp_table[11'h271] <= 9'h00e; exp_table[11'h272] <= 9'h00e; exp_table[11'h273] <= 9'h00e; exp_table[11'h274] <= 9'h00e; exp_table[11'h275] <= 9'h00e; exp_table[11'h276] <= 9'h00e; exp_table[11'h277] <= 9'h00e; exp_table[11'h278] <= 9'h00e; exp_table[11'h279] <= 9'h00e; exp_table[11'h27a] <= 9'h00e; exp_table[11'h27b] <= 9'h00e; exp_table[11'h27c] <= 9'h00d; exp_table[11'h27d] <= 9'h00d; exp_table[11'h27e] <= 9'h00d; exp_table[11'h27f] <= 9'h00d;
    exp_table[11'h280] <= 9'h00d; exp_table[11'h281] <= 9'h00d; exp_table[11'h282] <= 9'h00d; exp_table[11'h283] <= 9'h00d; exp_table[11'h284] <= 9'h00d; exp_table[11'h285] <= 9'h00d; exp_table[11'h286] <= 9'h00d; exp_table[11'h287] <= 9'h00d; exp_table[11'h288] <= 9'h00d; exp_table[11'h289] <= 9'h00d; exp_table[11'h28a] <= 9'h00c; exp_table[11'h28b] <= 9'h00c; exp_table[11'h28c] <= 9'h00c; exp_table[11'h28d] <= 9'h00c; exp_table[11'h28e] <= 9'h00c; exp_table[11'h28f] <= 9'h00c;
    exp_table[11'h290] <= 9'h00c; exp_table[11'h291] <= 9'h00c; exp_table[11'h292] <= 9'h00c; exp_table[11'h293] <= 9'h00c; exp_table[11'h294] <= 9'h00c; exp_table[11'h295] <= 9'h00c; exp_table[11'h296] <= 9'h00c; exp_table[11'h297] <= 9'h00c; exp_table[11'h298] <= 9'h00b; exp_table[11'h299] <= 9'h00b; exp_table[11'h29a] <= 9'h00b; exp_table[11'h29b] <= 9'h00b; exp_table[11'h29c] <= 9'h00b; exp_table[11'h29d] <= 9'h00b; exp_table[11'h29e] <= 9'h00b; exp_table[11'h29f] <= 9'h00b;
    exp_table[11'h2a0] <= 9'h00b; exp_table[11'h2a1] <= 9'h00b; exp_table[11'h2a2] <= 9'h00b; exp_table[11'h2a3] <= 9'h00b; exp_table[11'h2a4] <= 9'h00b; exp_table[11'h2a5] <= 9'h00b; exp_table[11'h2a6] <= 9'h00b; exp_table[11'h2a7] <= 9'h00a; exp_table[11'h2a8] <= 9'h00a; exp_table[11'h2a9] <= 9'h00a; exp_table[11'h2aa] <= 9'h00a; exp_table[11'h2ab] <= 9'h00a; exp_table[11'h2ac] <= 9'h00a; exp_table[11'h2ad] <= 9'h00a; exp_table[11'h2ae] <= 9'h00a; exp_table[11'h2af] <= 9'h00a;
    exp_table[11'h2b0] <= 9'h00a; exp_table[11'h2b1] <= 9'h00a; exp_table[11'h2b2] <= 9'h00a; exp_table[11'h2b3] <= 9'h00a; exp_table[11'h2b4] <= 9'h00a; exp_table[11'h2b5] <= 9'h00a; exp_table[11'h2b6] <= 9'h00a; exp_table[11'h2b7] <= 9'h00a; exp_table[11'h2b8] <= 9'h009; exp_table[11'h2b9] <= 9'h009; exp_table[11'h2ba] <= 9'h009; exp_table[11'h2bb] <= 9'h009; exp_table[11'h2bc] <= 9'h009; exp_table[11'h2bd] <= 9'h009; exp_table[11'h2be] <= 9'h009; exp_table[11'h2bf] <= 9'h009;
    exp_table[11'h2c0] <= 9'h009; exp_table[11'h2c1] <= 9'h009; exp_table[11'h2c2] <= 9'h009; exp_table[11'h2c3] <= 9'h009; exp_table[11'h2c4] <= 9'h009; exp_table[11'h2c5] <= 9'h009; exp_table[11'h2c6] <= 9'h009; exp_table[11'h2c7] <= 9'h009; exp_table[11'h2c8] <= 9'h009; exp_table[11'h2c9] <= 9'h009; exp_table[11'h2ca] <= 9'h009; exp_table[11'h2cb] <= 9'h008; exp_table[11'h2cc] <= 9'h008; exp_table[11'h2cd] <= 9'h008; exp_table[11'h2ce] <= 9'h008; exp_table[11'h2cf] <= 9'h008;
    exp_table[11'h2d0] <= 9'h008; exp_table[11'h2d1] <= 9'h008; exp_table[11'h2d2] <= 9'h008; exp_table[11'h2d3] <= 9'h008; exp_table[11'h2d4] <= 9'h008; exp_table[11'h2d5] <= 9'h008; exp_table[11'h2d6] <= 9'h008; exp_table[11'h2d7] <= 9'h008; exp_table[11'h2d8] <= 9'h008; exp_table[11'h2d9] <= 9'h008; exp_table[11'h2da] <= 9'h008; exp_table[11'h2db] <= 9'h008; exp_table[11'h2dc] <= 9'h008; exp_table[11'h2dd] <= 9'h008; exp_table[11'h2de] <= 9'h008; exp_table[11'h2df] <= 9'h007;
    exp_table[11'h2e0] <= 9'h007; exp_table[11'h2e1] <= 9'h007; exp_table[11'h2e2] <= 9'h007; exp_table[11'h2e3] <= 9'h007; exp_table[11'h2e4] <= 9'h007; exp_table[11'h2e5] <= 9'h007; exp_table[11'h2e6] <= 9'h007; exp_table[11'h2e7] <= 9'h007; exp_table[11'h2e8] <= 9'h007; exp_table[11'h2e9] <= 9'h007; exp_table[11'h2ea] <= 9'h007; exp_table[11'h2eb] <= 9'h007; exp_table[11'h2ec] <= 9'h007; exp_table[11'h2ed] <= 9'h007; exp_table[11'h2ee] <= 9'h007; exp_table[11'h2ef] <= 9'h007;
    exp_table[11'h2f0] <= 9'h007; exp_table[11'h2f1] <= 9'h007; exp_table[11'h2f2] <= 9'h007; exp_table[11'h2f3] <= 9'h007; exp_table[11'h2f4] <= 9'h007; exp_table[11'h2f5] <= 9'h007; exp_table[11'h2f6] <= 9'h007; exp_table[11'h2f7] <= 9'h006; exp_table[11'h2f8] <= 9'h006; exp_table[11'h2f9] <= 9'h006; exp_table[11'h2fa] <= 9'h006; exp_table[11'h2fb] <= 9'h006; exp_table[11'h2fc] <= 9'h006; exp_table[11'h2fd] <= 9'h006; exp_table[11'h2fe] <= 9'h006; exp_table[11'h2ff] <= 9'h006;
    exp_table[11'h300] <= 9'h006; exp_table[11'h301] <= 9'h006; exp_table[11'h302] <= 9'h006; exp_table[11'h303] <= 9'h006; exp_table[11'h304] <= 9'h006; exp_table[11'h305] <= 9'h006; exp_table[11'h306] <= 9'h006; exp_table[11'h307] <= 9'h006; exp_table[11'h308] <= 9'h006; exp_table[11'h309] <= 9'h006; exp_table[11'h30a] <= 9'h006; exp_table[11'h30b] <= 9'h006; exp_table[11'h30c] <= 9'h006; exp_table[11'h30d] <= 9'h006; exp_table[11'h30e] <= 9'h006; exp_table[11'h30f] <= 9'h006;
    exp_table[11'h310] <= 9'h006; exp_table[11'h311] <= 9'h006; exp_table[11'h312] <= 9'h005; exp_table[11'h313] <= 9'h005; exp_table[11'h314] <= 9'h005; exp_table[11'h315] <= 9'h005; exp_table[11'h316] <= 9'h005; exp_table[11'h317] <= 9'h005; exp_table[11'h318] <= 9'h005; exp_table[11'h319] <= 9'h005; exp_table[11'h31a] <= 9'h005; exp_table[11'h31b] <= 9'h005; exp_table[11'h31c] <= 9'h005; exp_table[11'h31d] <= 9'h005; exp_table[11'h31e] <= 9'h005; exp_table[11'h31f] <= 9'h005;
    exp_table[11'h320] <= 9'h005; exp_table[11'h321] <= 9'h005; exp_table[11'h322] <= 9'h005; exp_table[11'h323] <= 9'h005; exp_table[11'h324] <= 9'h005; exp_table[11'h325] <= 9'h005; exp_table[11'h326] <= 9'h005; exp_table[11'h327] <= 9'h005; exp_table[11'h328] <= 9'h005; exp_table[11'h329] <= 9'h005; exp_table[11'h32a] <= 9'h005; exp_table[11'h32b] <= 9'h005; exp_table[11'h32c] <= 9'h005; exp_table[11'h32d] <= 9'h005; exp_table[11'h32e] <= 9'h005; exp_table[11'h32f] <= 9'h005;
    exp_table[11'h330] <= 9'h005; exp_table[11'h331] <= 9'h005; exp_table[11'h332] <= 9'h004; exp_table[11'h333] <= 9'h004; exp_table[11'h334] <= 9'h004; exp_table[11'h335] <= 9'h004; exp_table[11'h336] <= 9'h004; exp_table[11'h337] <= 9'h004; exp_table[11'h338] <= 9'h004; exp_table[11'h339] <= 9'h004; exp_table[11'h33a] <= 9'h004; exp_table[11'h33b] <= 9'h004; exp_table[11'h33c] <= 9'h004; exp_table[11'h33d] <= 9'h004; exp_table[11'h33e] <= 9'h004; exp_table[11'h33f] <= 9'h004;
    exp_table[11'h340] <= 9'h004; exp_table[11'h341] <= 9'h004; exp_table[11'h342] <= 9'h004; exp_table[11'h343] <= 9'h004; exp_table[11'h344] <= 9'h004; exp_table[11'h345] <= 9'h004; exp_table[11'h346] <= 9'h004; exp_table[11'h347] <= 9'h004; exp_table[11'h348] <= 9'h004; exp_table[11'h349] <= 9'h004; exp_table[11'h34a] <= 9'h004; exp_table[11'h34b] <= 9'h004; exp_table[11'h34c] <= 9'h004; exp_table[11'h34d] <= 9'h004; exp_table[11'h34e] <= 9'h004; exp_table[11'h34f] <= 9'h004;
    exp_table[11'h350] <= 9'h004; exp_table[11'h351] <= 9'h004; exp_table[11'h352] <= 9'h004; exp_table[11'h353] <= 9'h004; exp_table[11'h354] <= 9'h004; exp_table[11'h355] <= 9'h004; exp_table[11'h356] <= 9'h004; exp_table[11'h357] <= 9'h004; exp_table[11'h358] <= 9'h004; exp_table[11'h359] <= 9'h004; exp_table[11'h35a] <= 9'h003; exp_table[11'h35b] <= 9'h003; exp_table[11'h35c] <= 9'h003; exp_table[11'h35d] <= 9'h003; exp_table[11'h35e] <= 9'h003; exp_table[11'h35f] <= 9'h003;
    exp_table[11'h360] <= 9'h003; exp_table[11'h361] <= 9'h003; exp_table[11'h362] <= 9'h003; exp_table[11'h363] <= 9'h003; exp_table[11'h364] <= 9'h003; exp_table[11'h365] <= 9'h003; exp_table[11'h366] <= 9'h003; exp_table[11'h367] <= 9'h003; exp_table[11'h368] <= 9'h003; exp_table[11'h369] <= 9'h003; exp_table[11'h36a] <= 9'h003; exp_table[11'h36b] <= 9'h003; exp_table[11'h36c] <= 9'h003; exp_table[11'h36d] <= 9'h003; exp_table[11'h36e] <= 9'h003; exp_table[11'h36f] <= 9'h003;
    exp_table[11'h370] <= 9'h003; exp_table[11'h371] <= 9'h003; exp_table[11'h372] <= 9'h003; exp_table[11'h373] <= 9'h003; exp_table[11'h374] <= 9'h003; exp_table[11'h375] <= 9'h003; exp_table[11'h376] <= 9'h003; exp_table[11'h377] <= 9'h003; exp_table[11'h378] <= 9'h003; exp_table[11'h379] <= 9'h003; exp_table[11'h37a] <= 9'h003; exp_table[11'h37b] <= 9'h003; exp_table[11'h37c] <= 9'h003; exp_table[11'h37d] <= 9'h003; exp_table[11'h37e] <= 9'h003; exp_table[11'h37f] <= 9'h003;
    exp_table[11'h380] <= 9'h003; exp_table[11'h381] <= 9'h003; exp_table[11'h382] <= 9'h003; exp_table[11'h383] <= 9'h003; exp_table[11'h384] <= 9'h003; exp_table[11'h385] <= 9'h003; exp_table[11'h386] <= 9'h003; exp_table[11'h387] <= 9'h003; exp_table[11'h388] <= 9'h003; exp_table[11'h389] <= 9'h003; exp_table[11'h38a] <= 9'h003; exp_table[11'h38b] <= 9'h003; exp_table[11'h38c] <= 9'h003; exp_table[11'h38d] <= 9'h002; exp_table[11'h38e] <= 9'h002; exp_table[11'h38f] <= 9'h002;
    exp_table[11'h390] <= 9'h002; exp_table[11'h391] <= 9'h002; exp_table[11'h392] <= 9'h002; exp_table[11'h393] <= 9'h002; exp_table[11'h394] <= 9'h002; exp_table[11'h395] <= 9'h002; exp_table[11'h396] <= 9'h002; exp_table[11'h397] <= 9'h002; exp_table[11'h398] <= 9'h002; exp_table[11'h399] <= 9'h002; exp_table[11'h39a] <= 9'h002; exp_table[11'h39b] <= 9'h002; exp_table[11'h39c] <= 9'h002; exp_table[11'h39d] <= 9'h002; exp_table[11'h39e] <= 9'h002; exp_table[11'h39f] <= 9'h002;
    exp_table[11'h3a0] <= 9'h002; exp_table[11'h3a1] <= 9'h002; exp_table[11'h3a2] <= 9'h002; exp_table[11'h3a3] <= 9'h002; exp_table[11'h3a4] <= 9'h002; exp_table[11'h3a5] <= 9'h002; exp_table[11'h3a6] <= 9'h002; exp_table[11'h3a7] <= 9'h002; exp_table[11'h3a8] <= 9'h002; exp_table[11'h3a9] <= 9'h002; exp_table[11'h3aa] <= 9'h002; exp_table[11'h3ab] <= 9'h002; exp_table[11'h3ac] <= 9'h002; exp_table[11'h3ad] <= 9'h002; exp_table[11'h3ae] <= 9'h002; exp_table[11'h3af] <= 9'h002;
    exp_table[11'h3b0] <= 9'h002; exp_table[11'h3b1] <= 9'h002; exp_table[11'h3b2] <= 9'h002; exp_table[11'h3b3] <= 9'h002; exp_table[11'h3b4] <= 9'h002; exp_table[11'h3b5] <= 9'h002; exp_table[11'h3b6] <= 9'h002; exp_table[11'h3b7] <= 9'h002; exp_table[11'h3b8] <= 9'h002; exp_table[11'h3b9] <= 9'h002; exp_table[11'h3ba] <= 9'h002; exp_table[11'h3bb] <= 9'h002; exp_table[11'h3bc] <= 9'h002; exp_table[11'h3bd] <= 9'h002; exp_table[11'h3be] <= 9'h002; exp_table[11'h3bf] <= 9'h002;
    exp_table[11'h3c0] <= 9'h002; exp_table[11'h3c1] <= 9'h002; exp_table[11'h3c2] <= 9'h002; exp_table[11'h3c3] <= 9'h002; exp_table[11'h3c4] <= 9'h002; exp_table[11'h3c5] <= 9'h002; exp_table[11'h3c6] <= 9'h002; exp_table[11'h3c7] <= 9'h002; exp_table[11'h3c8] <= 9'h002; exp_table[11'h3c9] <= 9'h002; exp_table[11'h3ca] <= 9'h002; exp_table[11'h3cb] <= 9'h002; exp_table[11'h3cc] <= 9'h002; exp_table[11'h3cd] <= 9'h002; exp_table[11'h3ce] <= 9'h002; exp_table[11'h3cf] <= 9'h002;
    exp_table[11'h3d0] <= 9'h002; exp_table[11'h3d1] <= 9'h002; exp_table[11'h3d2] <= 9'h002; exp_table[11'h3d3] <= 9'h002; exp_table[11'h3d4] <= 9'h001; exp_table[11'h3d5] <= 9'h001; exp_table[11'h3d6] <= 9'h001; exp_table[11'h3d7] <= 9'h001; exp_table[11'h3d8] <= 9'h001; exp_table[11'h3d9] <= 9'h001; exp_table[11'h3da] <= 9'h001; exp_table[11'h3db] <= 9'h001; exp_table[11'h3dc] <= 9'h001; exp_table[11'h3dd] <= 9'h001; exp_table[11'h3de] <= 9'h001; exp_table[11'h3df] <= 9'h001;
    exp_table[11'h3e0] <= 9'h001; exp_table[11'h3e1] <= 9'h001; exp_table[11'h3e2] <= 9'h001; exp_table[11'h3e3] <= 9'h001; exp_table[11'h3e4] <= 9'h001; exp_table[11'h3e5] <= 9'h001; exp_table[11'h3e6] <= 9'h001; exp_table[11'h3e7] <= 9'h001; exp_table[11'h3e8] <= 9'h001; exp_table[11'h3e9] <= 9'h001; exp_table[11'h3ea] <= 9'h001; exp_table[11'h3eb] <= 9'h001; exp_table[11'h3ec] <= 9'h001; exp_table[11'h3ed] <= 9'h001; exp_table[11'h3ee] <= 9'h001; exp_table[11'h3ef] <= 9'h001;
    exp_table[11'h3f0] <= 9'h001; exp_table[11'h3f1] <= 9'h001; exp_table[11'h3f2] <= 9'h001; exp_table[11'h3f3] <= 9'h001; exp_table[11'h3f4] <= 9'h001; exp_table[11'h3f5] <= 9'h001; exp_table[11'h3f6] <= 9'h001; exp_table[11'h3f7] <= 9'h001; exp_table[11'h3f8] <= 9'h001; exp_table[11'h3f9] <= 9'h001; exp_table[11'h3fa] <= 9'h001; exp_table[11'h3fb] <= 9'h001; exp_table[11'h3fc] <= 9'h001; exp_table[11'h3fd] <= 9'h001; exp_table[11'h3fe] <= 9'h001; exp_table[11'h3ff] <= 9'h001;
end

always @ (posedge clk) begin
    value <= ((addr[10] == 0) && (addr[11] == 0)) ? exp_table[addr] : 0;
end

endmodule
